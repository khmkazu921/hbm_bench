`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/21/2020 01:48:45 PM
// Design Name: 
// Module Name: combine
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module combine
  #(
    parameter int MOD_NUM = 32,
    parameter int COUNT_NUM = 34,
    parameter int DATA_WIDTH = 256
    )
    (
     input SYS_CLK0_N,
     input SYS_CLK0_P
     );
    
    wire   clk_450;
    wire   aresetn_450;

    AXI3 axi3  [0:MOD_NUM-1]();
    Monitor mon[0:MOD_NUM-1]();

    reg [39:0] count;
    wire       iswrite;
    wire       isread = ~iswrite;
    wire [3:0] state;
    wire random;
    wire [3:0] len;
    wire [4:0] select_port;
    
    // always_ff @(posedge clk_450) begin
    //     if(aresetn_450 == 0) 
    //       count <= 0;            
    //     else 
    //       count <= ~count[39] ? count + 1 : count;
    // end
    
    generate
        for(genvar i = 0; i < MOD_NUM; i = i + 1) begin: GenFloattester_0
            assign mon[i].isread = isread;
            assign mon[i].iswrite = iswrite;
            assign mon[i].state = state;
            assign mon[i].random = random;
            assign mon[i].len = len;
            //assign mon[i].select_port = select_port;
            float_tester_top #(.DATA_WIDTH(DATA_WIDTH), .MOD_RANK(i), .PORT_RANK(i)) float_tester_top_0
              ( .aclk(clk_450), .aresetn(aresetn_450), .axi3(axi3[i]), .mon(mon[i]) );  
        end        
    endgenerate

    wire clk_100;
    wire locked;
    wire trigger;
    wire resetn;

    clk_wiz_0 clk_wiz_0_inst
      (
       .clk_in1_n(SYS_CLK0_N),
       .clk_in1_p(SYS_CLK0_P),
       .clk_100(clk_100),
       .clk_450(clk_450),
       .locked(locked)
       );

    user_reset user_reset_inst
      (
       .clk(clk_450),
       .trigger(trigger),
       .mig_rstn(resetn)
       );

    proc_sys_reset_0 proc_sys_reset_450
      (
       .slowest_sync_clk(clk_450),
       .ext_reset_in(1),
       .aux_reset_in(resetn),
       .mb_debug_sys_rst(0),
       .dcm_locked(locked),
       .peripheral_aresetn(aresetn_450)
       );
    
//    ila_0 ila_0_inst
//      (
//       .clk(clk_450),
//       .probe0 (mon[0 ].awaddr),
//       );

    vio_0 vio_0_inst
      (
       .clk(clk_450),
       .probe_out0(trigger),
       .probe_out1(state),
       .probe_out2(random),
       .probe_out3(iswrite),
       .probe_out4 (len),
       .probe_out5 (mon[0].select_port),
       .probe_out6 (mon[1].select_port),
       .probe_out7 (mon[2].select_port),
       .probe_out8 (mon[3].select_port),
       .probe_out9 (mon[4].select_port),
       .probe_out10(mon[5].select_port),
       .probe_out11(mon[6].select_port),
       .probe_out12(mon[7].select_port),
       .probe_out13(mon[8].select_port),
       .probe_out14(mon[9].select_port),
       .probe_out15(mon[10].select_port),
       .probe_out16(mon[11].select_port),
       .probe_out17(mon[12].select_port),
       .probe_out18(mon[13].select_port),
       .probe_out19(mon[14].select_port),
       .probe_out20(mon[15].select_port),
       .probe_out21(mon[16].select_port),
       .probe_out22(mon[17].select_port),
       .probe_out23(mon[18].select_port),
       .probe_out24(mon[19].select_port),
       .probe_out25(mon[20].select_port),
       .probe_out26(mon[21].select_port),
       .probe_out27(mon[22].select_port),
       .probe_out28(mon[23].select_port),
       .probe_out29(mon[24].select_port),
       .probe_out30(mon[25].select_port),
       .probe_out31(mon[26].select_port),
       .probe_out32(mon[27].select_port),
       .probe_out33(mon[28].select_port),
       .probe_out34(mon[29].select_port),
       .probe_out35(mon[30].select_port),
       .probe_out36(mon[31].select_port)
       );
       
    vio_1 vio_1_inst
      (
       .clk(clk_450),
       .probe_out0(mon[0].reset),
       .probe_out1(mon[1].reset),
       .probe_out2(mon[2].reset),
       .probe_out3(mon[3].reset),
       .probe_out4(mon[4].reset),
       .probe_out5(mon[5].reset),
       .probe_out6(mon[6].reset),
       .probe_out7(mon[7].reset),
       .probe_out8(mon[8].reset),
       .probe_out9(mon[9].reset),
       .probe_out10(mon[10].reset),
       .probe_out11(mon[11].reset),
       .probe_out12(mon[12].reset),
       .probe_out13(mon[13].reset),
       .probe_out14(mon[14].reset),
       .probe_out15(mon[15].reset),
       .probe_out16(mon[16].reset),
       .probe_out17(mon[17].reset),
       .probe_out18(mon[18].reset),
       .probe_out19(mon[19].reset),
       .probe_out20(mon[20].reset),
       .probe_out21(mon[21].reset),
       .probe_out22(mon[22].reset),
       .probe_out23(mon[23].reset),
       .probe_out24(mon[24].reset),
       .probe_out25(mon[25].reset),
       .probe_out26(mon[26].reset),
       .probe_out27(mon[27].reset),
       .probe_out28(mon[28].reset),
       .probe_out29(mon[29].reset),
       .probe_out30(mon[30].reset),
       .probe_out31(mon[31].reset)
       );
       
    hbm_0 hbm_0_inst 
     (
      .APB_0_PCLK         (clk_100            ),
      .APB_0_PRESET_N     (resetn             ),
      .apb_complete_0     (                   ),
      .DRAM_0_STAT_CATTRIP(                   ),
      .DRAM_0_STAT_TEMP   (                   ),
      .HBM_REF_CLK_0      (clk_450            ),
      .APB_1_PCLK         (clk_100            ),
      .APB_1_PRESET_N     (resetn             ),
      .apb_complete_1     (                   ),
      .DRAM_1_STAT_CATTRIP(                   ),
      .DRAM_1_STAT_TEMP   (                   ),
      .HBM_REF_CLK_1      (clk_450            ),
      .AXI_00_ACLK        (clk_450            ),
      .AXI_00_ARESET_N    (aresetn_450        ),
      .AXI_00_ARADDR      (axi3[0].araddr     ),
      .AXI_00_ARBURST     (axi3[0].arburst    ),
      .AXI_00_ARID        (axi3[0].arid       ),
      .AXI_00_ARLEN       (axi3[0].arlen      ),
      .AXI_00_ARSIZE      (axi3[0].arsize     ),
      .AXI_00_ARVALID     (axi3[0].arvalid    ),
      .AXI_00_AWADDR      (axi3[0].awaddr     ),
      .AXI_00_AWBURST     (axi3[0].awburst    ),
      .AXI_00_AWID        (axi3[0].awid       ),
      .AXI_00_AWLEN       (axi3[0].awlen      ),
      .AXI_00_AWSIZE      (axi3[0].awsize     ),
      .AXI_00_AWVALID     (axi3[0].awvalid    ),
      .AXI_00_RREADY      (axi3[0].rready     ),
      .AXI_00_BREADY      (axi3[0].bready     ),
      .AXI_00_WDATA       (axi3[0].wdata      ),
      .AXI_00_WLAST       (axi3[0].wlast      ),
      .AXI_00_WSTRB       (axi3[0].wstrb      ),
      .AXI_00_WDATA_PARITY(                   ), 
      .AXI_00_WVALID      (axi3[0].wvalid     ),
      .AXI_00_ARREADY     (axi3[0].arready    ),
      .AXI_00_AWREADY     (axi3[0].awready    ),
      .AXI_00_RDATA_PARITY(                   ), 
      .AXI_00_RDATA       (axi3[0].rdata      ),
      .AXI_00_RID         (axi3[0].rid        ),
      .AXI_00_RLAST       (axi3[0].rlast      ),
      .AXI_00_RRESP       (axi3[0].rresp      ),
      .AXI_00_RVALID      (axi3[0].rvalid     ),
      .AXI_00_WREADY      (axi3[0].wready     ),
      .AXI_00_BID         (axi3[0].bid        ),
      .AXI_00_BRESP       (axi3[0].bresp      ),
      .AXI_00_BVALID      (axi3[0].bvalid     ),
      .AXI_01_ACLK        (clk_450            ),
      .AXI_01_ARESET_N    (aresetn_450        ),
      .AXI_01_ARADDR      (axi3[1].araddr     ),
      .AXI_01_ARBURST     (axi3[1].arburst    ),
      .AXI_01_ARID        (axi3[1].arid       ),
      .AXI_01_ARLEN       (axi3[1].arlen      ),
      .AXI_01_ARSIZE      (axi3[1].arsize     ),
      .AXI_01_ARVALID     (axi3[1].arvalid    ),
      .AXI_01_AWADDR      (axi3[1].awaddr     ),
      .AXI_01_AWBURST     (axi3[1].awburst    ),
      .AXI_01_AWID        (axi3[1].awid       ),
      .AXI_01_AWLEN       (axi3[1].awlen      ),
      .AXI_01_AWSIZE      (axi3[1].awsize     ),
      .AXI_01_AWVALID     (axi3[1].awvalid    ),
      .AXI_01_RREADY      (axi3[1].rready     ),
      .AXI_01_BREADY      (axi3[1].bready     ),
      .AXI_01_WDATA       (axi3[1].wdata      ),
      .AXI_01_WLAST       (axi3[1].wlast      ),
      .AXI_01_WSTRB       (axi3[1].wstrb      ),
      .AXI_01_WDATA_PARITY(                   ), 
      .AXI_01_WVALID      (axi3[1].wvalid     ),
      .AXI_01_ARREADY     (axi3[1].arready    ),
      .AXI_01_AWREADY     (axi3[1].awready    ),
      .AXI_01_RDATA_PARITY(                   ), 
      .AXI_01_RDATA       (axi3[1].rdata      ),
      .AXI_01_RID         (axi3[1].rid        ),
      .AXI_01_RLAST       (axi3[1].rlast      ),
      .AXI_01_RRESP       (axi3[1].rresp      ),
      .AXI_01_RVALID      (axi3[1].rvalid     ),
      .AXI_01_WREADY      (axi3[1].wready     ),
      .AXI_01_BID         (axi3[1].bid        ),
      .AXI_01_BRESP       (axi3[1].bresp      ),
      .AXI_01_BVALID      (axi3[1].bvalid     ),
      .AXI_02_ACLK        (clk_450            ),
      .AXI_02_ARESET_N    (aresetn_450        ),
      .AXI_02_ARADDR      (axi3[2].araddr     ),
      .AXI_02_ARBURST     (axi3[2].arburst    ),
      .AXI_02_ARID        (axi3[2].arid       ),
      .AXI_02_ARLEN       (axi3[2].arlen      ),
      .AXI_02_ARSIZE      (axi3[2].arsize     ),
      .AXI_02_ARVALID     (axi3[2].arvalid    ),
      .AXI_02_AWADDR      (axi3[2].awaddr     ),
      .AXI_02_AWBURST     (axi3[2].awburst    ),
      .AXI_02_AWID        (axi3[2].awid       ),
      .AXI_02_AWLEN       (axi3[2].awlen      ),
      .AXI_02_AWSIZE      (axi3[2].awsize     ),
      .AXI_02_AWVALID     (axi3[2].awvalid    ),
      .AXI_02_RREADY      (axi3[2].rready     ),
      .AXI_02_BREADY      (axi3[2].bready     ),
      .AXI_02_WDATA       (axi3[2].wdata      ),
      .AXI_02_WLAST       (axi3[2].wlast      ),
      .AXI_02_WSTRB       (axi3[2].wstrb      ),
      .AXI_02_WDATA_PARITY(                   ),
      .AXI_02_WVALID      (axi3[2].wvalid     ),
      .AXI_02_ARREADY     (axi3[2].arready    ),
      .AXI_02_AWREADY     (axi3[2].awready    ),
      .AXI_02_RDATA_PARITY(                   ),
      .AXI_02_RDATA       (axi3[2].rdata      ),
      .AXI_02_RID         (axi3[2].rid        ),
      .AXI_02_RLAST       (axi3[2].rlast      ),
      .AXI_02_RRESP       (axi3[2].rresp      ),
      .AXI_02_RVALID      (axi3[2].rvalid     ),
      .AXI_02_WREADY      (axi3[2].wready     ),
      .AXI_02_BID         (axi3[2].bid        ),
      .AXI_02_BRESP       (axi3[2].bresp      ),
      .AXI_02_BVALID      (axi3[2].bvalid     ),
      .AXI_03_ACLK        (clk_450            ),
      .AXI_03_ARESET_N    (aresetn_450        ),
      .AXI_03_ARADDR      (axi3[3].araddr     ),
      .AXI_03_ARBURST     (axi3[3].arburst    ),
      .AXI_03_ARID        (axi3[3].arid       ),
      .AXI_03_ARLEN       (axi3[3].arlen      ),
      .AXI_03_ARSIZE      (axi3[3].arsize     ),
      .AXI_03_ARVALID     (axi3[3].arvalid    ),
      .AXI_03_AWADDR      (axi3[3].awaddr     ),
      .AXI_03_AWBURST     (axi3[3].awburst    ),
      .AXI_03_AWID        (axi3[3].awid       ),
      .AXI_03_AWLEN       (axi3[3].awlen      ),
      .AXI_03_AWSIZE      (axi3[3].awsize     ),
      .AXI_03_AWVALID     (axi3[3].awvalid    ),
      .AXI_03_RREADY      (axi3[3].rready     ),
      .AXI_03_BREADY      (axi3[3].bready     ),
      .AXI_03_WDATA       (axi3[3].wdata      ),
      .AXI_03_WLAST       (axi3[3].wlast      ),
      .AXI_03_WSTRB       (axi3[3].wstrb      ),
      .AXI_03_WDATA_PARITY(                   ),
      .AXI_03_WVALID      (axi3[3].wvalid     ),
      .AXI_03_ARREADY     (axi3[3].arready    ),
      .AXI_03_AWREADY     (axi3[3].awready    ),
      .AXI_03_RDATA_PARITY(                   ),
      .AXI_03_RDATA       (axi3[3].rdata      ),
      .AXI_03_RID         (axi3[3].rid        ),
      .AXI_03_RLAST       (axi3[3].rlast      ),
      .AXI_03_RRESP       (axi3[3].rresp      ),
      .AXI_03_RVALID      (axi3[3].rvalid     ),
      .AXI_03_WREADY      (axi3[3].wready     ),
      .AXI_03_BID         (axi3[3].bid        ),
      .AXI_03_BRESP       (axi3[3].bresp      ),
      .AXI_03_BVALID      (axi3[3].bvalid     ),
      .AXI_04_ACLK        (clk_450            ),
      .AXI_04_ARESET_N    (aresetn_450        ),
      .AXI_04_ARADDR      (axi3[4].araddr     ),
      .AXI_04_ARBURST     (axi3[4].arburst    ),
      .AXI_04_ARID        (axi3[4].arid       ),
      .AXI_04_ARLEN       (axi3[4].arlen      ),
      .AXI_04_ARSIZE      (axi3[4].arsize     ),
      .AXI_04_ARVALID     (axi3[4].arvalid    ),
      .AXI_04_AWADDR      (axi3[4].awaddr     ),
      .AXI_04_AWBURST     (axi3[4].awburst    ),
      .AXI_04_AWID        (axi3[4].awid       ),
      .AXI_04_AWLEN       (axi3[4].awlen      ),
      .AXI_04_AWSIZE      (axi3[4].awsize     ),
      .AXI_04_AWVALID     (axi3[4].awvalid    ),
      .AXI_04_RREADY      (axi3[4].rready     ),
      .AXI_04_BREADY      (axi3[4].bready     ),
      .AXI_04_WDATA       (axi3[4].wdata      ),
      .AXI_04_WLAST       (axi3[4].wlast      ),
      .AXI_04_WSTRB       (axi3[4].wstrb      ),
      .AXI_04_WDATA_PARITY(                   ),
      .AXI_04_WVALID      (axi3[4].wvalid     ),
      .AXI_04_ARREADY     (axi3[4].arready    ),
      .AXI_04_AWREADY     (axi3[4].awready    ),
      .AXI_04_RDATA_PARITY(                   ),
      .AXI_04_RDATA       (axi3[4].rdata      ),
      .AXI_04_RID         (axi3[4].rid        ),
      .AXI_04_RLAST       (axi3[4].rlast      ),
      .AXI_04_RRESP       (axi3[4].rresp      ),
      .AXI_04_RVALID      (axi3[4].rvalid     ),
      .AXI_04_WREADY      (axi3[4].wready     ),
      .AXI_04_BID         (axi3[4].bid        ),
      .AXI_04_BRESP       (axi3[4].bresp      ),
      .AXI_04_BVALID      (axi3[4].bvalid     ),
      .AXI_05_ACLK        (clk_450            ),
      .AXI_05_ARESET_N    (aresetn_450        ),
      .AXI_05_ARADDR      (axi3[5].araddr     ),
      .AXI_05_ARBURST     (axi3[5].arburst    ),
      .AXI_05_ARID        (axi3[5].arid       ),
      .AXI_05_ARLEN       (axi3[5].arlen      ),
      .AXI_05_ARSIZE      (axi3[5].arsize     ),
      .AXI_05_ARVALID     (axi3[5].arvalid    ),
      .AXI_05_AWADDR      (axi3[5].awaddr     ),
      .AXI_05_AWBURST     (axi3[5].awburst    ),
      .AXI_05_AWID        (axi3[5].awid       ),
      .AXI_05_AWLEN       (axi3[5].awlen      ),
      .AXI_05_AWSIZE      (axi3[5].awsize     ),
      .AXI_05_AWVALID     (axi3[5].awvalid    ),
      .AXI_05_RREADY      (axi3[5].rready     ),
      .AXI_05_BREADY      (axi3[5].bready     ),
      .AXI_05_WDATA       (axi3[5].wdata      ),
      .AXI_05_WLAST       (axi3[5].wlast      ),
      .AXI_05_WSTRB       (axi3[5].wstrb      ),
      .AXI_05_WDATA_PARITY(                   ),
      .AXI_05_WVALID      (axi3[5].wvalid     ),
      .AXI_05_ARREADY     (axi3[5].arready    ),
      .AXI_05_AWREADY     (axi3[5].awready    ),
      .AXI_05_RDATA_PARITY(                   ),
      .AXI_05_RDATA       (axi3[5].rdata      ),
      .AXI_05_RID         (axi3[5].rid        ),
      .AXI_05_RLAST       (axi3[5].rlast      ),
      .AXI_05_RRESP       (axi3[5].rresp      ),
      .AXI_05_RVALID      (axi3[5].rvalid     ),
      .AXI_05_WREADY      (axi3[5].wready     ),
      .AXI_05_BID         (axi3[5].bid        ),
      .AXI_05_BRESP       (axi3[5].bresp      ),
      .AXI_05_BVALID      (axi3[5].bvalid     ),
      .AXI_06_ACLK        (clk_450            ),
      .AXI_06_ARESET_N    (aresetn_450        ),
      .AXI_06_ARADDR      (axi3[6].araddr     ),
      .AXI_06_ARBURST     (axi3[6].arburst    ),
      .AXI_06_ARID        (axi3[6].arid       ),
      .AXI_06_ARLEN       (axi3[6].arlen      ),
      .AXI_06_ARSIZE      (axi3[6].arsize     ),
      .AXI_06_ARVALID     (axi3[6].arvalid    ),
      .AXI_06_AWADDR      (axi3[6].awaddr     ),
      .AXI_06_AWBURST     (axi3[6].awburst    ),
      .AXI_06_AWID        (axi3[6].awid       ),
      .AXI_06_AWLEN       (axi3[6].awlen      ),
      .AXI_06_AWSIZE      (axi3[6].awsize     ),
      .AXI_06_AWVALID     (axi3[6].awvalid    ),
      .AXI_06_RREADY      (axi3[6].rready     ),
      .AXI_06_BREADY      (axi3[6].bready     ),
      .AXI_06_WDATA       (axi3[6].wdata      ),
      .AXI_06_WLAST       (axi3[6].wlast      ),
      .AXI_06_WSTRB       (axi3[6].wstrb      ),
      .AXI_06_WDATA_PARITY(                   ),
      .AXI_06_WVALID      (axi3[6].wvalid     ),
      .AXI_06_ARREADY     (axi3[6].arready    ),
      .AXI_06_AWREADY     (axi3[6].awready    ),
      .AXI_06_RDATA_PARITY(                   ),
      .AXI_06_RDATA       (axi3[6].rdata      ),
      .AXI_06_RID         (axi3[6].rid        ),
      .AXI_06_RLAST       (axi3[6].rlast      ),
      .AXI_06_RRESP       (axi3[6].rresp      ),
      .AXI_06_RVALID      (axi3[6].rvalid     ),
      .AXI_06_WREADY      (axi3[6].wready     ),
      .AXI_06_BID         (axi3[6].bid        ),
      .AXI_06_BRESP       (axi3[6].bresp      ),
      .AXI_06_BVALID      (axi3[6].bvalid     ),
      .AXI_07_ACLK        (clk_450            ),
      .AXI_07_ARESET_N    (aresetn_450        ),
      .AXI_07_ARADDR      (axi3[7].araddr     ),
      .AXI_07_ARBURST     (axi3[7].arburst    ),
      .AXI_07_ARID        (axi3[7].arid       ),
      .AXI_07_ARLEN       (axi3[7].arlen      ),
      .AXI_07_ARSIZE      (axi3[7].arsize     ),
      .AXI_07_ARVALID     (axi3[7].arvalid    ),
      .AXI_07_AWADDR      (axi3[7].awaddr     ),
      .AXI_07_AWBURST     (axi3[7].awburst    ),
      .AXI_07_AWID        (axi3[7].awid       ),
      .AXI_07_AWLEN       (axi3[7].awlen      ),
      .AXI_07_AWSIZE      (axi3[7].awsize     ),
      .AXI_07_AWVALID     (axi3[7].awvalid    ),
      .AXI_07_RREADY      (axi3[7].rready     ),
      .AXI_07_BREADY      (axi3[7].bready     ),
      .AXI_07_WDATA       (axi3[7].wdata      ),
      .AXI_07_WLAST       (axi3[7].wlast      ),
      .AXI_07_WSTRB       (axi3[7].wstrb      ),
      .AXI_07_WDATA_PARITY(                   ),
      .AXI_07_WVALID      (axi3[7].wvalid     ),
      .AXI_07_ARREADY     (axi3[7].arready    ),
      .AXI_07_AWREADY     (axi3[7].awready    ),
      .AXI_07_RDATA_PARITY(                   ),
      .AXI_07_RDATA       (axi3[7].rdata      ),
      .AXI_07_RID         (axi3[7].rid        ),
      .AXI_07_RLAST       (axi3[7].rlast      ),
      .AXI_07_RRESP       (axi3[7].rresp      ),
      .AXI_07_RVALID      (axi3[7].rvalid     ),
      .AXI_07_WREADY      (axi3[7].wready     ),
      .AXI_07_BID         (axi3[7].bid        ),
      .AXI_07_BRESP       (axi3[7].bresp      ),
      .AXI_07_BVALID      (axi3[7].bvalid     ),
      .AXI_08_ACLK        (clk_450            ),
      .AXI_08_ARESET_N    (aresetn_450        ),
      .AXI_08_ARADDR      (axi3[8].araddr     ),
      .AXI_08_ARBURST     (axi3[8].arburst    ),
      .AXI_08_ARID        (axi3[8].arid       ),
      .AXI_08_ARLEN       (axi3[8].arlen      ),
      .AXI_08_ARSIZE      (axi3[8].arsize     ),
      .AXI_08_ARVALID     (axi3[8].arvalid    ),
      .AXI_08_AWADDR      (axi3[8].awaddr     ),
      .AXI_08_AWBURST     (axi3[8].awburst    ),
      .AXI_08_AWID        (axi3[8].awid       ),
      .AXI_08_AWLEN       (axi3[8].awlen      ),
      .AXI_08_AWSIZE      (axi3[8].awsize     ),
      .AXI_08_AWVALID     (axi3[8].awvalid    ),
      .AXI_08_RREADY      (axi3[8].rready     ),
      .AXI_08_BREADY      (axi3[8].bready     ),
      .AXI_08_WDATA       (axi3[8].wdata      ),
      .AXI_08_WLAST       (axi3[8].wlast      ),
      .AXI_08_WSTRB       (axi3[8].wstrb      ),
      .AXI_08_WDATA_PARITY(                   ),
      .AXI_08_WVALID      (axi3[8].wvalid     ),
      .AXI_08_ARREADY     (axi3[8].arready    ),
      .AXI_08_AWREADY     (axi3[8].awready    ),
      .AXI_08_RDATA_PARITY(                   ),
      .AXI_08_RDATA       (axi3[8].rdata      ),
      .AXI_08_RID         (axi3[8].rid        ),
      .AXI_08_RLAST       (axi3[8].rlast      ),
      .AXI_08_RRESP       (axi3[8].rresp      ),
      .AXI_08_RVALID      (axi3[8].rvalid     ),
      .AXI_08_WREADY      (axi3[8].wready     ),
      .AXI_08_BID         (axi3[8].bid        ),
      .AXI_08_BRESP       (axi3[8].bresp      ),
      .AXI_08_BVALID      (axi3[8].bvalid     ),
      .AXI_09_ACLK        (clk_450            ),
      .AXI_09_ARESET_N    (aresetn_450        ),
      .AXI_09_ARADDR      (axi3[9].araddr     ),
      .AXI_09_ARBURST     (axi3[9].arburst    ),
      .AXI_09_ARID        (axi3[9].arid       ),
      .AXI_09_ARLEN       (axi3[9].arlen      ),
      .AXI_09_ARSIZE      (axi3[9].arsize     ),
      .AXI_09_ARVALID     (axi3[9].arvalid    ),
      .AXI_09_AWADDR      (axi3[9].awaddr     ),
      .AXI_09_AWBURST     (axi3[9].awburst    ),
      .AXI_09_AWID        (axi3[9].awid       ),
      .AXI_09_AWLEN       (axi3[9].awlen      ),
      .AXI_09_AWSIZE      (axi3[9].awsize     ),
      .AXI_09_AWVALID     (axi3[9].awvalid    ),
      .AXI_09_RREADY      (axi3[9].rready     ),
      .AXI_09_BREADY      (axi3[9].bready     ),
      .AXI_09_WDATA       (axi3[9].wdata      ),
      .AXI_09_WLAST       (axi3[9].wlast      ),
      .AXI_09_WSTRB       (axi3[9].wstrb      ),
      .AXI_09_WDATA_PARITY(                   ),
      .AXI_09_WVALID      (axi3[9].wvalid     ),
      .AXI_09_ARREADY     (axi3[9].arready    ),
      .AXI_09_AWREADY     (axi3[9].awready    ),
      .AXI_09_RDATA_PARITY(                   ),
      .AXI_09_RDATA       (axi3[9].rdata      ),
      .AXI_09_RID         (axi3[9].rid        ),
      .AXI_09_RLAST       (axi3[9].rlast      ),
      .AXI_09_RRESP       (axi3[9].rresp      ),
      .AXI_09_RVALID      (axi3[9].rvalid     ),
      .AXI_09_WREADY      (axi3[9].wready     ),
      .AXI_09_BID         (axi3[9].bid        ),
      .AXI_09_BRESP       (axi3[9].bresp      ),
      .AXI_09_BVALID      (axi3[9].bvalid     ),
      .AXI_10_ACLK        (clk_450            ),
      .AXI_10_ARESET_N    (aresetn_450        ),
      .AXI_10_ARADDR      (axi3[10].araddr    ),
      .AXI_10_ARBURST     (axi3[10].arburst   ),
      .AXI_10_ARID        (axi3[10].arid      ),
      .AXI_10_ARLEN       (axi3[10].arlen     ),
      .AXI_10_ARSIZE      (axi3[10].arsize    ),
      .AXI_10_ARVALID     (axi3[10].arvalid   ),
      .AXI_10_AWADDR      (axi3[10].awaddr    ),
      .AXI_10_AWBURST     (axi3[10].awburst   ),
      .AXI_10_AWID        (axi3[10].awid      ),
      .AXI_10_AWLEN       (axi3[10].awlen     ),
      .AXI_10_AWSIZE      (axi3[10].awsize    ),
      .AXI_10_AWVALID     (axi3[10].awvalid   ),
      .AXI_10_RREADY      (axi3[10].rready    ),
      .AXI_10_BREADY      (axi3[10].bready    ),
      .AXI_10_WDATA       (axi3[10].wdata     ),
      .AXI_10_WLAST       (axi3[10].wlast     ),
      .AXI_10_WSTRB       (axi3[10].wstrb     ),
      .AXI_10_WDATA_PARITY(                   ),
      .AXI_10_WVALID      (axi3[10].wvalid    ),
      .AXI_10_ARREADY     (axi3[10].arready   ),
      .AXI_10_AWREADY     (axi3[10].awready   ),
      .AXI_10_RDATA_PARITY(                   ),
      .AXI_10_RDATA       (axi3[10].rdata     ),
      .AXI_10_RID         (axi3[10].rid       ),
      .AXI_10_RLAST       (axi3[10].rlast     ),
      .AXI_10_RRESP       (axi3[10].rresp     ),
      .AXI_10_RVALID      (axi3[10].rvalid    ),
      .AXI_10_WREADY      (axi3[10].wready    ),
      .AXI_10_BID         (axi3[10].bid       ),
      .AXI_10_BRESP       (axi3[10].bresp     ),
      .AXI_10_BVALID      (axi3[10].bvalid    ),
      .AXI_11_ACLK        (clk_450            ),
      .AXI_11_ARESET_N    (aresetn_450        ),
      .AXI_11_ARADDR      (axi3[11].araddr    ),
      .AXI_11_ARBURST     (axi3[11].arburst   ),
      .AXI_11_ARID        (axi3[11].arid      ),
      .AXI_11_ARLEN       (axi3[11].arlen     ),
      .AXI_11_ARSIZE      (axi3[11].arsize    ),
      .AXI_11_ARVALID     (axi3[11].arvalid   ),
      .AXI_11_AWADDR      (axi3[11].awaddr    ),
      .AXI_11_AWBURST     (axi3[11].awburst   ),
      .AXI_11_AWID        (axi3[11].awid      ),
      .AXI_11_AWLEN       (axi3[11].awlen     ),
      .AXI_11_AWSIZE      (axi3[11].awsize    ),
      .AXI_11_AWVALID     (axi3[11].awvalid   ),
      .AXI_11_RREADY      (axi3[11].rready    ),
      .AXI_11_BREADY      (axi3[11].bready    ),
      .AXI_11_WDATA       (axi3[11].wdata     ),
      .AXI_11_WLAST       (axi3[11].wlast     ),
      .AXI_11_WSTRB       (axi3[11].wstrb     ),
      .AXI_11_WDATA_PARITY(                   ),
      .AXI_11_WVALID      (axi3[11].wvalid    ),
      .AXI_11_ARREADY     (axi3[11].arready   ),
      .AXI_11_AWREADY     (axi3[11].awready   ),
      .AXI_11_RDATA_PARITY(                   ),
      .AXI_11_RDATA       (axi3[11].rdata     ),
      .AXI_11_RID         (axi3[11].rid       ),
      .AXI_11_RLAST       (axi3[11].rlast     ),
      .AXI_11_RRESP       (axi3[11].rresp     ),
      .AXI_11_RVALID      (axi3[11].rvalid    ),
      .AXI_11_WREADY      (axi3[11].wready    ),
      .AXI_11_BID         (axi3[11].bid       ),
      .AXI_11_BRESP       (axi3[11].bresp     ),
      .AXI_11_BVALID      (axi3[11].bvalid    ),
      .AXI_12_ACLK        (clk_450            ),
      .AXI_12_ARESET_N    (aresetn_450        ),
      .AXI_12_ARADDR      (axi3[12].araddr    ),
      .AXI_12_ARBURST     (axi3[12].arburst   ),
      .AXI_12_ARID        (axi3[12].arid      ),
      .AXI_12_ARLEN       (axi3[12].arlen     ),
      .AXI_12_ARSIZE      (axi3[12].arsize    ),
      .AXI_12_ARVALID     (axi3[12].arvalid   ),
      .AXI_12_AWADDR      (axi3[12].awaddr    ),
      .AXI_12_AWBURST     (axi3[12].awburst   ),
      .AXI_12_AWID        (axi3[12].awid      ),
      .AXI_12_AWLEN       (axi3[12].awlen     ),
      .AXI_12_AWSIZE      (axi3[12].awsize    ),
      .AXI_12_AWVALID     (axi3[12].awvalid   ),
      .AXI_12_RREADY      (axi3[12].rready    ),
      .AXI_12_BREADY      (axi3[12].bready    ),
      .AXI_12_WDATA       (axi3[12].wdata     ),
      .AXI_12_WLAST       (axi3[12].wlast     ),
      .AXI_12_WSTRB       (axi3[12].wstrb     ),
      .AXI_12_WDATA_PARITY(                   ),
      .AXI_12_WVALID      (axi3[12].wvalid    ),
      .AXI_12_ARREADY     (axi3[12].arready   ),
      .AXI_12_AWREADY     (axi3[12].awready   ),
      .AXI_12_RDATA_PARITY(                   ),
      .AXI_12_RDATA       (axi3[12].rdata     ),
      .AXI_12_RID         (axi3[12].rid       ),
      .AXI_12_RLAST       (axi3[12].rlast     ),
      .AXI_12_RRESP       (axi3[12].rresp     ),
      .AXI_12_RVALID      (axi3[12].rvalid    ),
      .AXI_12_WREADY      (axi3[12].wready    ),
      .AXI_12_BID         (axi3[12].bid       ),
      .AXI_12_BRESP       (axi3[12].bresp     ),
      .AXI_12_BVALID      (axi3[12].bvalid    ),
      .AXI_13_ACLK        (clk_450            ),
      .AXI_13_ARESET_N    (aresetn_450        ),
      .AXI_13_ARADDR      (axi3[13].araddr    ),
      .AXI_13_ARBURST     (axi3[13].arburst   ),
      .AXI_13_ARID        (axi3[13].arid      ),
      .AXI_13_ARLEN       (axi3[13].arlen     ),
      .AXI_13_ARSIZE      (axi3[13].arsize    ),
      .AXI_13_ARVALID     (axi3[13].arvalid   ),
      .AXI_13_AWADDR      (axi3[13].awaddr    ),
      .AXI_13_AWBURST     (axi3[13].awburst   ),
      .AXI_13_AWID        (axi3[13].awid      ),
      .AXI_13_AWLEN       (axi3[13].awlen     ),
      .AXI_13_AWSIZE      (axi3[13].awsize    ),
      .AXI_13_AWVALID     (axi3[13].awvalid   ),
      .AXI_13_RREADY      (axi3[13].rready    ),
      .AXI_13_BREADY      (axi3[13].bready    ),
      .AXI_13_WDATA       (axi3[13].wdata     ),
      .AXI_13_WLAST       (axi3[13].wlast     ),
      .AXI_13_WSTRB       (axi3[13].wstrb     ),
      .AXI_13_WDATA_PARITY(                   ),
      .AXI_13_WVALID      (axi3[13].wvalid    ),
      .AXI_13_ARREADY     (axi3[13].arready   ),
      .AXI_13_AWREADY     (axi3[13].awready   ),
      .AXI_13_RDATA_PARITY(                   ),
      .AXI_13_RDATA       (axi3[13].rdata     ),
      .AXI_13_RID         (axi3[13].rid       ),
      .AXI_13_RLAST       (axi3[13].rlast     ),
      .AXI_13_RRESP       (axi3[13].rresp     ),
      .AXI_13_RVALID      (axi3[13].rvalid    ),
      .AXI_13_WREADY      (axi3[13].wready    ),
      .AXI_13_BID         (axi3[13].bid       ),
      .AXI_13_BRESP       (axi3[13].bresp     ),
      .AXI_13_BVALID      (axi3[13].bvalid    ),
      .AXI_14_ACLK        (clk_450            ),
      .AXI_14_ARESET_N    (aresetn_450        ),
      .AXI_14_ARADDR      (axi3[14].araddr    ),
      .AXI_14_ARBURST     (axi3[14].arburst   ),
      .AXI_14_ARID        (axi3[14].arid      ),
      .AXI_14_ARLEN       (axi3[14].arlen     ),
      .AXI_14_ARSIZE      (axi3[14].arsize    ),
      .AXI_14_ARVALID     (axi3[14].arvalid   ),
      .AXI_14_AWADDR      (axi3[14].awaddr    ),
      .AXI_14_AWBURST     (axi3[14].awburst   ),
      .AXI_14_AWID        (axi3[14].awid      ),
      .AXI_14_AWLEN       (axi3[14].awlen     ),
      .AXI_14_AWSIZE      (axi3[14].awsize    ),
      .AXI_14_AWVALID     (axi3[14].awvalid   ),
      .AXI_14_RREADY      (axi3[14].rready    ),
      .AXI_14_BREADY      (axi3[14].bready    ),
      .AXI_14_WDATA       (axi3[14].wdata     ),
      .AXI_14_WLAST       (axi3[14].wlast     ),
      .AXI_14_WSTRB       (axi3[14].wstrb     ),
      .AXI_14_WDATA_PARITY(                   ),
      .AXI_14_WVALID      (axi3[14].wvalid    ),
      .AXI_14_ARREADY     (axi3[14].arready   ),
      .AXI_14_AWREADY     (axi3[14].awready   ),
      .AXI_14_RDATA_PARITY(                   ),
      .AXI_14_RDATA       (axi3[14].rdata     ),
      .AXI_14_RID         (axi3[14].rid       ),
      .AXI_14_RLAST       (axi3[14].rlast     ),
      .AXI_14_RRESP       (axi3[14].rresp     ),
      .AXI_14_RVALID      (axi3[14].rvalid    ),
      .AXI_14_WREADY      (axi3[14].wready    ),
      .AXI_14_BID         (axi3[14].bid       ),
      .AXI_14_BRESP       (axi3[14].bresp     ),
      .AXI_14_BVALID      (axi3[14].bvalid    ),
      .AXI_15_ACLK        (clk_450            ),
      .AXI_15_ARESET_N    (aresetn_450        ),
      .AXI_15_ARADDR      (axi3[15].araddr    ),
      .AXI_15_ARBURST     (axi3[15].arburst   ),
      .AXI_15_ARID        (axi3[15].arid      ),
      .AXI_15_ARLEN       (axi3[15].arlen     ),
      .AXI_15_ARSIZE      (axi3[15].arsize    ),
      .AXI_15_ARVALID     (axi3[15].arvalid   ),
      .AXI_15_AWADDR      (axi3[15].awaddr    ),
      .AXI_15_AWBURST     (axi3[15].awburst   ),
      .AXI_15_AWID        (axi3[15].awid      ),
      .AXI_15_AWLEN       (axi3[15].awlen     ),
      .AXI_15_AWSIZE      (axi3[15].awsize    ),
      .AXI_15_AWVALID     (axi3[15].awvalid   ),
      .AXI_15_RREADY      (axi3[15].rready    ),
      .AXI_15_BREADY      (axi3[15].bready    ),
      .AXI_15_WDATA       (axi3[15].wdata     ),
      .AXI_15_WLAST       (axi3[15].wlast     ),
      .AXI_15_WSTRB       (axi3[15].wstrb     ),
      .AXI_15_WDATA_PARITY(                   ),
      .AXI_15_WVALID      (axi3[15].wvalid    ),
      .AXI_15_ARREADY     (axi3[15].arready   ),
      .AXI_15_AWREADY     (axi3[15].awready   ),
      .AXI_15_RDATA_PARITY(                   ),
      .AXI_15_RDATA       (axi3[15].rdata     ),
      .AXI_15_RID         (axi3[15].rid       ),
      .AXI_15_RLAST       (axi3[15].rlast     ),
      .AXI_15_RRESP       (axi3[15].rresp     ),
      .AXI_15_RVALID      (axi3[15].rvalid    ),
      .AXI_15_WREADY      (axi3[15].wready    ),
      .AXI_15_BID         (axi3[15].bid       ),
      .AXI_15_BRESP       (axi3[15].bresp     ),
      .AXI_15_BVALID      (axi3[15].bvalid    ),
      .AXI_16_ACLK        (clk_450            ),
      .AXI_16_ARESET_N    (aresetn_450        ),
      .AXI_16_ARADDR      (axi3[16].araddr    ),
      .AXI_16_ARBURST     (axi3[16].arburst   ),
      .AXI_16_ARID        (axi3[16].arid      ),
      .AXI_16_ARLEN       (axi3[16].arlen     ),
      .AXI_16_ARSIZE      (axi3[16].arsize    ),
      .AXI_16_ARVALID     (axi3[16].arvalid   ),
      .AXI_16_AWADDR      (axi3[16].awaddr    ),
      .AXI_16_AWBURST     (axi3[16].awburst   ),
      .AXI_16_AWID        (axi3[16].awid      ),
      .AXI_16_AWLEN       (axi3[16].awlen     ),
      .AXI_16_AWSIZE      (axi3[16].awsize    ),
      .AXI_16_AWVALID     (axi3[16].awvalid   ),
      .AXI_16_RREADY      (axi3[16].rready    ),
      .AXI_16_BREADY      (axi3[16].bready    ),
      .AXI_16_WDATA       (axi3[16].wdata     ),
      .AXI_16_WLAST       (axi3[16].wlast     ),
      .AXI_16_WSTRB       (axi3[16].wstrb     ),
      .AXI_16_WDATA_PARITY(                   ),
      .AXI_16_WVALID      (axi3[16].wvalid    ),
      .AXI_16_ARREADY     (axi3[16].arready   ),
      .AXI_16_AWREADY     (axi3[16].awready   ),
      .AXI_16_RDATA_PARITY(                   ),
      .AXI_16_RDATA       (axi3[16].rdata     ),
      .AXI_16_RID         (axi3[16].rid       ),
      .AXI_16_RLAST       (axi3[16].rlast     ),
      .AXI_16_RRESP       (axi3[16].rresp     ),
      .AXI_16_RVALID      (axi3[16].rvalid    ),
      .AXI_16_WREADY      (axi3[16].wready    ),
      .AXI_16_BID         (axi3[16].bid       ),
      .AXI_16_BRESP       (axi3[16].bresp     ),
      .AXI_16_BVALID      (axi3[16].bvalid    ),
      .AXI_17_ACLK        (clk_450            ),
      .AXI_17_ARESET_N    (aresetn_450        ),
      .AXI_17_ARADDR      (axi3[17].araddr    ),
      .AXI_17_ARBURST     (axi3[17].arburst   ),
      .AXI_17_ARID        (axi3[17].arid      ),
      .AXI_17_ARLEN       (axi3[17].arlen     ),
      .AXI_17_ARSIZE      (axi3[17].arsize    ),
      .AXI_17_ARVALID     (axi3[17].arvalid   ),
      .AXI_17_AWADDR      (axi3[17].awaddr    ),
      .AXI_17_AWBURST     (axi3[17].awburst   ),
      .AXI_17_AWID        (axi3[17].awid      ),
      .AXI_17_AWLEN       (axi3[17].awlen     ),
      .AXI_17_AWSIZE      (axi3[17].awsize    ),
      .AXI_17_AWVALID     (axi3[17].awvalid   ),
      .AXI_17_RREADY      (axi3[17].rready    ),
      .AXI_17_BREADY      (axi3[17].bready    ),
      .AXI_17_WDATA       (axi3[17].wdata     ),
      .AXI_17_WLAST       (axi3[17].wlast     ),
      .AXI_17_WSTRB       (axi3[17].wstrb     ),
      .AXI_17_WDATA_PARITY(                   ),
      .AXI_17_WVALID      (axi3[17].wvalid    ),
      .AXI_17_ARREADY     (axi3[17].arready   ),
      .AXI_17_AWREADY     (axi3[17].awready   ),
      .AXI_17_RDATA_PARITY(                   ),
      .AXI_17_RDATA       (axi3[17].rdata     ),
      .AXI_17_RID         (axi3[17].rid       ),
      .AXI_17_RLAST       (axi3[17].rlast     ),
      .AXI_17_RRESP       (axi3[17].rresp     ),
      .AXI_17_RVALID      (axi3[17].rvalid    ),
      .AXI_17_WREADY      (axi3[17].wready    ),
      .AXI_17_BID         (axi3[17].bid       ),
      .AXI_17_BRESP       (axi3[17].bresp     ),
      .AXI_17_BVALID      (axi3[17].bvalid    ),
      .AXI_18_ACLK        (clk_450            ),
      .AXI_18_ARESET_N    (aresetn_450        ),
      .AXI_18_ARADDR      (axi3[18].araddr    ),
      .AXI_18_ARBURST     (axi3[18].arburst   ),
      .AXI_18_ARID        (axi3[18].arid      ),
      .AXI_18_ARLEN       (axi3[18].arlen     ),
      .AXI_18_ARSIZE      (axi3[18].arsize    ),
      .AXI_18_ARVALID     (axi3[18].arvalid   ),
      .AXI_18_AWADDR      (axi3[18].awaddr    ),
      .AXI_18_AWBURST     (axi3[18].awburst   ),
      .AXI_18_AWID        (axi3[18].awid      ),
      .AXI_18_AWLEN       (axi3[18].awlen     ),
      .AXI_18_AWSIZE      (axi3[18].awsize    ),
      .AXI_18_AWVALID     (axi3[18].awvalid   ),
      .AXI_18_RREADY      (axi3[18].rready    ),
      .AXI_18_BREADY      (axi3[18].bready    ),
      .AXI_18_WDATA       (axi3[18].wdata     ),
      .AXI_18_WLAST       (axi3[18].wlast     ),
      .AXI_18_WSTRB       (axi3[18].wstrb     ),
      .AXI_18_WDATA_PARITY(                   ),
      .AXI_18_WVALID      (axi3[18].wvalid    ),
      .AXI_18_ARREADY     (axi3[18].arready   ),
      .AXI_18_AWREADY     (axi3[18].awready   ),
      .AXI_18_RDATA_PARITY(                   ),
      .AXI_18_RDATA       (axi3[18].rdata     ),
      .AXI_18_RID         (axi3[18].rid       ),
      .AXI_18_RLAST       (axi3[18].rlast     ),
      .AXI_18_RRESP       (axi3[18].rresp     ),
      .AXI_18_RVALID      (axi3[18].rvalid    ),
      .AXI_18_WREADY      (axi3[18].wready    ),
      .AXI_18_BID         (axi3[18].bid       ),
      .AXI_18_BRESP       (axi3[18].bresp     ),
      .AXI_18_BVALID      (axi3[18].bvalid    ),
      .AXI_19_ACLK        (clk_450            ),
      .AXI_19_ARESET_N    (aresetn_450        ),
      .AXI_19_ARADDR      (axi3[19].araddr    ),
      .AXI_19_ARBURST     (axi3[19].arburst   ),
      .AXI_19_ARID        (axi3[19].arid      ),
      .AXI_19_ARLEN       (axi3[19].arlen     ),
      .AXI_19_ARSIZE      (axi3[19].arsize    ),
      .AXI_19_ARVALID     (axi3[19].arvalid   ),
      .AXI_19_AWADDR      (axi3[19].awaddr    ),
      .AXI_19_AWBURST     (axi3[19].awburst   ),
      .AXI_19_AWID        (axi3[19].awid      ),
      .AXI_19_AWLEN       (axi3[19].awlen     ),
      .AXI_19_AWSIZE      (axi3[19].awsize    ),
      .AXI_19_AWVALID     (axi3[19].awvalid   ),
      .AXI_19_RREADY      (axi3[19].rready    ),
      .AXI_19_BREADY      (axi3[19].bready    ),
      .AXI_19_WDATA       (axi3[19].wdata     ),
      .AXI_19_WLAST       (axi3[19].wlast     ),
      .AXI_19_WSTRB       (axi3[19].wstrb     ),
      .AXI_19_WDATA_PARITY(                   ),
      .AXI_19_WVALID      (axi3[19].wvalid    ),
      .AXI_19_ARREADY     (axi3[19].arready   ),
      .AXI_19_AWREADY     (axi3[19].awready   ),
      .AXI_19_RDATA_PARITY(                   ),
      .AXI_19_RDATA       (axi3[19].rdata     ),
      .AXI_19_RID         (axi3[19].rid       ),
      .AXI_19_RLAST       (axi3[19].rlast     ),
      .AXI_19_RRESP       (axi3[19].rresp     ),
      .AXI_19_RVALID      (axi3[19].rvalid    ),
      .AXI_19_WREADY      (axi3[19].wready    ),
      .AXI_19_BID         (axi3[19].bid       ),
      .AXI_19_BRESP       (axi3[19].bresp     ),
      .AXI_19_BVALID      (axi3[19].bvalid    ),
      .AXI_20_ACLK        (clk_450            ),
      .AXI_20_ARESET_N    (aresetn_450        ),
      .AXI_20_ARADDR      (axi3[20].araddr    ),
      .AXI_20_ARBURST     (axi3[20].arburst   ),
      .AXI_20_ARID        (axi3[20].arid      ),
      .AXI_20_ARLEN       (axi3[20].arlen     ),
      .AXI_20_ARSIZE      (axi3[20].arsize    ),
      .AXI_20_ARVALID     (axi3[20].arvalid   ),
      .AXI_20_AWADDR      (axi3[20].awaddr    ),
      .AXI_20_AWBURST     (axi3[20].awburst   ),
      .AXI_20_AWID        (axi3[20].awid      ),
      .AXI_20_AWLEN       (axi3[20].awlen     ),
      .AXI_20_AWSIZE      (axi3[20].awsize    ),
      .AXI_20_AWVALID     (axi3[20].awvalid   ),
      .AXI_20_RREADY      (axi3[20].rready    ),
      .AXI_20_BREADY      (axi3[20].bready    ),
      .AXI_20_WDATA       (axi3[20].wdata     ),
      .AXI_20_WLAST       (axi3[20].wlast     ),
      .AXI_20_WSTRB       (axi3[20].wstrb     ),
      .AXI_20_WDATA_PARITY(                   ),
      .AXI_20_WVALID      (axi3[20].wvalid    ),
      .AXI_20_ARREADY     (axi3[20].arready   ),
      .AXI_20_AWREADY     (axi3[20].awready   ),
      .AXI_20_RDATA_PARITY(                   ),
      .AXI_20_RDATA       (axi3[20].rdata     ),
      .AXI_20_RID         (axi3[20].rid       ),
      .AXI_20_RLAST       (axi3[20].rlast     ),
      .AXI_20_RRESP       (axi3[20].rresp     ),
      .AXI_20_RVALID      (axi3[20].rvalid    ),
      .AXI_20_WREADY      (axi3[20].wready    ),
      .AXI_20_BID         (axi3[20].bid       ),
      .AXI_20_BRESP       (axi3[20].bresp     ),
      .AXI_20_BVALID      (axi3[20].bvalid    ),
      .AXI_21_ACLK        (clk_450            ),
      .AXI_21_ARESET_N    (aresetn_450        ),
      .AXI_21_ARADDR      (axi3[21].araddr    ),
      .AXI_21_ARBURST     (axi3[21].arburst   ),
      .AXI_21_ARID        (axi3[21].arid      ),
      .AXI_21_ARLEN       (axi3[21].arlen     ),
      .AXI_21_ARSIZE      (axi3[21].arsize    ),
      .AXI_21_ARVALID     (axi3[21].arvalid   ),
      .AXI_21_AWADDR      (axi3[21].awaddr    ),
      .AXI_21_AWBURST     (axi3[21].awburst   ),
      .AXI_21_AWID        (axi3[21].awid      ),
      .AXI_21_AWLEN       (axi3[21].awlen     ),
      .AXI_21_AWSIZE      (axi3[21].awsize    ),
      .AXI_21_AWVALID     (axi3[21].awvalid   ),
      .AXI_21_RREADY      (axi3[21].rready    ),
      .AXI_21_BREADY      (axi3[21].bready    ),
      .AXI_21_WDATA       (axi3[21].wdata     ),
      .AXI_21_WLAST       (axi3[21].wlast     ),
      .AXI_21_WSTRB       (axi3[21].wstrb     ),
      .AXI_21_WDATA_PARITY(                   ),
      .AXI_21_WVALID      (axi3[21].wvalid    ),
      .AXI_21_ARREADY     (axi3[21].arready   ),
      .AXI_21_AWREADY     (axi3[21].awready   ),
      .AXI_21_RDATA_PARITY(                   ),
      .AXI_21_RDATA       (axi3[21].rdata     ),
      .AXI_21_RID         (axi3[21].rid       ),
      .AXI_21_RLAST       (axi3[21].rlast     ),
      .AXI_21_RRESP       (axi3[21].rresp     ),
      .AXI_21_RVALID      (axi3[21].rvalid    ),
      .AXI_21_WREADY      (axi3[21].wready    ),
      .AXI_21_BID         (axi3[21].bid       ),
      .AXI_21_BRESP       (axi3[21].bresp     ),
      .AXI_21_BVALID      (axi3[21].bvalid    ),
      .AXI_22_ACLK        (clk_450            ),
      .AXI_22_ARESET_N    (aresetn_450        ),
      .AXI_22_ARADDR      (axi3[22].araddr    ),
      .AXI_22_ARBURST     (axi3[22].arburst   ),
      .AXI_22_ARID        (axi3[22].arid      ),
      .AXI_22_ARLEN       (axi3[22].arlen     ),
      .AXI_22_ARSIZE      (axi3[22].arsize    ),
      .AXI_22_ARVALID     (axi3[22].arvalid   ),
      .AXI_22_AWADDR      (axi3[22].awaddr    ),
      .AXI_22_AWBURST     (axi3[22].awburst   ),
      .AXI_22_AWID        (axi3[22].awid      ),
      .AXI_22_AWLEN       (axi3[22].awlen     ),
      .AXI_22_AWSIZE      (axi3[22].awsize    ),
      .AXI_22_AWVALID     (axi3[22].awvalid   ),
      .AXI_22_RREADY      (axi3[22].rready    ),
      .AXI_22_BREADY      (axi3[22].bready    ),
      .AXI_22_WDATA       (axi3[22].wdata     ),
      .AXI_22_WLAST       (axi3[22].wlast     ),
      .AXI_22_WSTRB       (axi3[22].wstrb     ),
      .AXI_22_WDATA_PARITY(                   ),
      .AXI_22_WVALID      (axi3[22].wvalid    ),
      .AXI_22_ARREADY     (axi3[22].arready   ),
      .AXI_22_AWREADY     (axi3[22].awready   ),
      .AXI_22_RDATA_PARITY(                   ),
      .AXI_22_RDATA       (axi3[22].rdata     ),
      .AXI_22_RID         (axi3[22].rid       ),
      .AXI_22_RLAST       (axi3[22].rlast     ),
      .AXI_22_RRESP       (axi3[22].rresp     ),
      .AXI_22_RVALID      (axi3[22].rvalid    ),
      .AXI_22_WREADY      (axi3[22].wready    ),
      .AXI_22_BID         (axi3[22].bid       ),
      .AXI_22_BRESP       (axi3[22].bresp     ),
      .AXI_22_BVALID      (axi3[22].bvalid    ),
      .AXI_23_ACLK        (clk_450            ),
      .AXI_23_ARESET_N    (aresetn_450        ),
      .AXI_23_ARADDR      (axi3[23].araddr    ),
      .AXI_23_ARBURST     (axi3[23].arburst   ),
      .AXI_23_ARID        (axi3[23].arid      ),
      .AXI_23_ARLEN       (axi3[23].arlen     ),
      .AXI_23_ARSIZE      (axi3[23].arsize    ),
      .AXI_23_ARVALID     (axi3[23].arvalid   ),
      .AXI_23_AWADDR      (axi3[23].awaddr    ),
      .AXI_23_AWBURST     (axi3[23].awburst   ),
      .AXI_23_AWID        (axi3[23].awid      ),
      .AXI_23_AWLEN       (axi3[23].awlen     ),
      .AXI_23_AWSIZE      (axi3[23].awsize    ),
      .AXI_23_AWVALID     (axi3[23].awvalid   ),
      .AXI_23_RREADY      (axi3[23].rready    ),
      .AXI_23_BREADY      (axi3[23].bready    ),
      .AXI_23_WDATA       (axi3[23].wdata     ),
      .AXI_23_WLAST       (axi3[23].wlast     ),
      .AXI_23_WSTRB       (axi3[23].wstrb     ),
      .AXI_23_WDATA_PARITY(                   ),
      .AXI_23_WVALID      (axi3[23].wvalid    ),
      .AXI_23_ARREADY     (axi3[23].arready   ),
      .AXI_23_AWREADY     (axi3[23].awready   ),
      .AXI_23_RDATA_PARITY(                   ),
      .AXI_23_RDATA       (axi3[23].rdata     ),
      .AXI_23_RID         (axi3[23].rid       ),
      .AXI_23_RLAST       (axi3[23].rlast     ),
      .AXI_23_RRESP       (axi3[23].rresp     ),
      .AXI_23_RVALID      (axi3[23].rvalid    ),
      .AXI_23_WREADY      (axi3[23].wready    ),
      .AXI_23_BID         (axi3[23].bid       ),
      .AXI_23_BRESP       (axi3[23].bresp     ),
      .AXI_23_BVALID      (axi3[23].bvalid    ),
      .AXI_24_ACLK        (clk_450            ),
      .AXI_24_ARESET_N    (aresetn_450        ),
      .AXI_24_ARADDR      (axi3[24].araddr    ),
      .AXI_24_ARBURST     (axi3[24].arburst   ),
      .AXI_24_ARID        (axi3[24].arid      ),
      .AXI_24_ARLEN       (axi3[24].arlen     ),
      .AXI_24_ARSIZE      (axi3[24].arsize    ),
      .AXI_24_ARVALID     (axi3[24].arvalid   ),
      .AXI_24_AWADDR      (axi3[24].awaddr    ),
      .AXI_24_AWBURST     (axi3[24].awburst   ),
      .AXI_24_AWID        (axi3[24].awid      ),
      .AXI_24_AWLEN       (axi3[24].awlen     ),
      .AXI_24_AWSIZE      (axi3[24].awsize    ),
      .AXI_24_AWVALID     (axi3[24].awvalid   ),
      .AXI_24_RREADY      (axi3[24].rready    ),
      .AXI_24_BREADY      (axi3[24].bready    ),
      .AXI_24_WDATA       (axi3[24].wdata     ),
      .AXI_24_WLAST       (axi3[24].wlast     ),
      .AXI_24_WSTRB       (axi3[24].wstrb     ),
      .AXI_24_WDATA_PARITY(                   ),
      .AXI_24_WVALID      (axi3[24].wvalid    ),
      .AXI_24_ARREADY     (axi3[24].arready   ),
      .AXI_24_AWREADY     (axi3[24].awready   ),
      .AXI_24_RDATA_PARITY(                   ),
      .AXI_24_RDATA       (axi3[24].rdata     ),
      .AXI_24_RID         (axi3[24].rid       ),
      .AXI_24_RLAST       (axi3[24].rlast     ),
      .AXI_24_RRESP       (axi3[24].rresp     ),
      .AXI_24_RVALID      (axi3[24].rvalid    ),
      .AXI_24_WREADY      (axi3[24].wready    ),
      .AXI_24_BID         (axi3[24].bid       ),
      .AXI_24_BRESP       (axi3[24].bresp     ),
      .AXI_24_BVALID      (axi3[24].bvalid    ),
      .AXI_25_ACLK        (clk_450            ),
      .AXI_25_ARESET_N    (aresetn_450        ),
      .AXI_25_ARADDR      (axi3[25].araddr    ),
      .AXI_25_ARBURST     (axi3[25].arburst   ),
      .AXI_25_ARID        (axi3[25].arid      ),
      .AXI_25_ARLEN       (axi3[25].arlen     ),
      .AXI_25_ARSIZE      (axi3[25].arsize    ),
      .AXI_25_ARVALID     (axi3[25].arvalid   ),
      .AXI_25_AWADDR      (axi3[25].awaddr    ),
      .AXI_25_AWBURST     (axi3[25].awburst   ),
      .AXI_25_AWID        (axi3[25].awid      ),
      .AXI_25_AWLEN       (axi3[25].awlen     ),
      .AXI_25_AWSIZE      (axi3[25].awsize    ),
      .AXI_25_AWVALID     (axi3[25].awvalid   ),
      .AXI_25_RREADY      (axi3[25].rready    ),
      .AXI_25_BREADY      (axi3[25].bready    ),
      .AXI_25_WDATA       (axi3[25].wdata     ),
      .AXI_25_WLAST       (axi3[25].wlast     ),
      .AXI_25_WSTRB       (axi3[25].wstrb     ),
      .AXI_25_WDATA_PARITY(                   ),
      .AXI_25_WVALID      (axi3[25].wvalid    ),
      .AXI_25_ARREADY     (axi3[25].arready   ),
      .AXI_25_AWREADY     (axi3[25].awready   ),
      .AXI_25_RDATA_PARITY(                   ),
      .AXI_25_RDATA       (axi3[25].rdata     ),
      .AXI_25_RID         (axi3[25].rid       ),
      .AXI_25_RLAST       (axi3[25].rlast     ),
      .AXI_25_RRESP       (axi3[25].rresp     ),
      .AXI_25_RVALID      (axi3[25].rvalid    ),
      .AXI_25_WREADY      (axi3[25].wready    ),
      .AXI_25_BID         (axi3[25].bid       ),
      .AXI_25_BRESP       (axi3[25].bresp     ),
      .AXI_25_BVALID      (axi3[25].bvalid    ),
      .AXI_26_ACLK        (clk_450            ),
      .AXI_26_ARESET_N    (aresetn_450        ),
      .AXI_26_ARADDR      (axi3[26].araddr    ),
      .AXI_26_ARBURST     (axi3[26].arburst   ),
      .AXI_26_ARID        (axi3[26].arid      ),
      .AXI_26_ARLEN       (axi3[26].arlen     ),
      .AXI_26_ARSIZE      (axi3[26].arsize    ),
      .AXI_26_ARVALID     (axi3[26].arvalid   ),
      .AXI_26_AWADDR      (axi3[26].awaddr    ),
      .AXI_26_AWBURST     (axi3[26].awburst   ),
      .AXI_26_AWID        (axi3[26].awid      ),
      .AXI_26_AWLEN       (axi3[26].awlen     ),
      .AXI_26_AWSIZE      (axi3[26].awsize    ),
      .AXI_26_AWVALID     (axi3[26].awvalid   ),
      .AXI_26_RREADY      (axi3[26].rready    ),
      .AXI_26_BREADY      (axi3[26].bready    ),
      .AXI_26_WDATA       (axi3[26].wdata     ),
      .AXI_26_WLAST       (axi3[26].wlast     ),
      .AXI_26_WSTRB       (axi3[26].wstrb     ),
      .AXI_26_WDATA_PARITY(                   ),
      .AXI_26_WVALID      (axi3[26].wvalid    ),
      .AXI_26_ARREADY     (axi3[26].arready   ),
      .AXI_26_AWREADY     (axi3[26].awready   ),
      .AXI_26_RDATA_PARITY(                   ),
      .AXI_26_RDATA       (axi3[26].rdata     ),
      .AXI_26_RID         (axi3[26].rid       ),
      .AXI_26_RLAST       (axi3[26].rlast     ),
      .AXI_26_RRESP       (axi3[26].rresp     ),
      .AXI_26_RVALID      (axi3[26].rvalid    ),
      .AXI_26_WREADY      (axi3[26].wready    ),
      .AXI_26_BID         (axi3[26].bid       ),
      .AXI_26_BRESP       (axi3[26].bresp     ),
      .AXI_26_BVALID      (axi3[26].bvalid    ),
      .AXI_27_ACLK        (clk_450            ),
      .AXI_27_ARESET_N    (aresetn_450        ),
      .AXI_27_ARADDR      (axi3[27].araddr    ),
      .AXI_27_ARBURST     (axi3[27].arburst   ),
      .AXI_27_ARID        (axi3[27].arid      ),
      .AXI_27_ARLEN       (axi3[27].arlen     ),
      .AXI_27_ARSIZE      (axi3[27].arsize    ),
      .AXI_27_ARVALID     (axi3[27].arvalid   ),
      .AXI_27_AWADDR      (axi3[27].awaddr    ),
      .AXI_27_AWBURST     (axi3[27].awburst   ),
      .AXI_27_AWID        (axi3[27].awid      ),
      .AXI_27_AWLEN       (axi3[27].awlen     ),
      .AXI_27_AWSIZE      (axi3[27].awsize    ),
      .AXI_27_AWVALID     (axi3[27].awvalid   ),
      .AXI_27_RREADY      (axi3[27].rready    ),
      .AXI_27_BREADY      (axi3[27].bready    ),
      .AXI_27_WDATA       (axi3[27].wdata     ),
      .AXI_27_WLAST       (axi3[27].wlast     ),
      .AXI_27_WSTRB       (axi3[27].wstrb     ),
      .AXI_27_WDATA_PARITY(                   ),
      .AXI_27_WVALID      (axi3[27].wvalid    ),
      .AXI_27_ARREADY     (axi3[27].arready   ),
      .AXI_27_AWREADY     (axi3[27].awready   ),
      .AXI_27_RDATA_PARITY(                   ),
      .AXI_27_RDATA       (axi3[27].rdata     ),
      .AXI_27_RID         (axi3[27].rid       ),
      .AXI_27_RLAST       (axi3[27].rlast     ),
      .AXI_27_RRESP       (axi3[27].rresp     ),
      .AXI_27_RVALID      (axi3[27].rvalid    ),
      .AXI_27_WREADY      (axi3[27].wready    ),
      .AXI_27_BID         (axi3[27].bid       ),
      .AXI_27_BRESP       (axi3[27].bresp     ),
      .AXI_27_BVALID      (axi3[27].bvalid    ),
      .AXI_28_ACLK        (clk_450            ),
      .AXI_28_ARESET_N    (aresetn_450        ),
      .AXI_28_ARADDR      (axi3[28].araddr    ),
      .AXI_28_ARBURST     (axi3[28].arburst   ),
      .AXI_28_ARID        (axi3[28].arid      ),
      .AXI_28_ARLEN       (axi3[28].arlen     ),
      .AXI_28_ARSIZE      (axi3[28].arsize    ),
      .AXI_28_ARVALID     (axi3[28].arvalid   ),
      .AXI_28_AWADDR      (axi3[28].awaddr    ),
      .AXI_28_AWBURST     (axi3[28].awburst   ),
      .AXI_28_AWID        (axi3[28].awid      ),
      .AXI_28_AWLEN       (axi3[28].awlen     ),
      .AXI_28_AWSIZE      (axi3[28].awsize    ),
      .AXI_28_AWVALID     (axi3[28].awvalid   ),
      .AXI_28_RREADY      (axi3[28].rready    ),
      .AXI_28_BREADY      (axi3[28].bready    ),
      .AXI_28_WDATA       (axi3[28].wdata     ),
      .AXI_28_WLAST       (axi3[28].wlast     ),
      .AXI_28_WSTRB       (axi3[28].wstrb     ),
      .AXI_28_WDATA_PARITY(                   ),
      .AXI_28_WVALID      (axi3[28].wvalid    ),
      .AXI_28_ARREADY     (axi3[28].arready   ),
      .AXI_28_AWREADY     (axi3[28].awready   ),
      .AXI_28_RDATA_PARITY(                   ),
      .AXI_28_RDATA       (axi3[28].rdata     ),
      .AXI_28_RID         (axi3[28].rid       ),
      .AXI_28_RLAST       (axi3[28].rlast     ),
      .AXI_28_RRESP       (axi3[28].rresp     ),
      .AXI_28_RVALID      (axi3[28].rvalid    ),
      .AXI_28_WREADY      (axi3[28].wready    ),
      .AXI_28_BID         (axi3[28].bid       ),
      .AXI_28_BRESP       (axi3[28].bresp     ),
      .AXI_28_BVALID      (axi3[28].bvalid    ),
      .AXI_29_ACLK        (clk_450            ),
      .AXI_29_ARESET_N    (aresetn_450        ),
      .AXI_29_ARADDR      (axi3[29].araddr    ),
      .AXI_29_ARBURST     (axi3[29].arburst   ),
      .AXI_29_ARID        (axi3[29].arid      ),
      .AXI_29_ARLEN       (axi3[29].arlen     ),
      .AXI_29_ARSIZE      (axi3[29].arsize    ),
      .AXI_29_ARVALID     (axi3[29].arvalid   ),
      .AXI_29_AWADDR      (axi3[29].awaddr    ),
      .AXI_29_AWBURST     (axi3[29].awburst   ),
      .AXI_29_AWID        (axi3[29].awid      ),
      .AXI_29_AWLEN       (axi3[29].awlen     ),
      .AXI_29_AWSIZE      (axi3[29].awsize    ),
      .AXI_29_AWVALID     (axi3[29].awvalid   ),
      .AXI_29_RREADY      (axi3[29].rready    ),
      .AXI_29_BREADY      (axi3[29].bready    ),
      .AXI_29_WDATA       (axi3[29].wdata     ),
      .AXI_29_WLAST       (axi3[29].wlast     ),
      .AXI_29_WSTRB       (axi3[29].wstrb     ),
      .AXI_29_WDATA_PARITY(                   ),
      .AXI_29_WVALID      (axi3[29].wvalid    ),
      .AXI_29_ARREADY     (axi3[29].arready   ),
      .AXI_29_AWREADY     (axi3[29].awready   ),
      .AXI_29_RDATA_PARITY(                   ),
      .AXI_29_RDATA       (axi3[29].rdata     ),
      .AXI_29_RID         (axi3[29].rid       ),
      .AXI_29_RLAST       (axi3[29].rlast     ),
      .AXI_29_RRESP       (axi3[29].rresp     ),
      .AXI_29_RVALID      (axi3[29].rvalid    ),
      .AXI_29_WREADY      (axi3[29].wready    ),
      .AXI_29_BID         (axi3[29].bid       ),
      .AXI_29_BRESP       (axi3[29].bresp     ),
      .AXI_29_BVALID      (axi3[29].bvalid    ),
      .AXI_30_ACLK        (clk_450            ),
      .AXI_30_ARESET_N    (aresetn_450        ),
      .AXI_30_ARADDR      (axi3[30].araddr    ),
      .AXI_30_ARBURST     (axi3[30].arburst   ),
      .AXI_30_ARID        (axi3[30].arid      ),
      .AXI_30_ARLEN       (axi3[30].arlen     ),
      .AXI_30_ARSIZE      (axi3[30].arsize    ),
      .AXI_30_ARVALID     (axi3[30].arvalid   ),
      .AXI_30_AWADDR      (axi3[30].awaddr    ),
      .AXI_30_AWBURST     (axi3[30].awburst   ),
      .AXI_30_AWID        (axi3[30].awid      ),
      .AXI_30_AWLEN       (axi3[30].awlen     ),
      .AXI_30_AWSIZE      (axi3[30].awsize    ),
      .AXI_30_AWVALID     (axi3[30].awvalid   ),
      .AXI_30_RREADY      (axi3[30].rready    ),
      .AXI_30_BREADY      (axi3[30].bready    ),
      .AXI_30_WDATA       (axi3[30].wdata     ),
      .AXI_30_WLAST       (axi3[30].wlast     ),
      .AXI_30_WSTRB       (axi3[30].wstrb     ),
      .AXI_30_WDATA_PARITY(                   ),
      .AXI_30_WVALID      (axi3[30].wvalid    ),
      .AXI_30_ARREADY     (axi3[30].arready   ),
      .AXI_30_AWREADY     (axi3[30].awready   ),
      .AXI_30_RDATA_PARITY(                   ),
      .AXI_30_RDATA       (axi3[30].rdata     ),
      .AXI_30_RID         (axi3[30].rid       ),
      .AXI_30_RLAST       (axi3[30].rlast     ),
      .AXI_30_RRESP       (axi3[30].rresp     ),
      .AXI_30_RVALID      (axi3[30].rvalid    ),
      .AXI_30_WREADY      (axi3[30].wready    ),
      .AXI_30_BID         (axi3[30].bid       ),
      .AXI_30_BRESP       (axi3[30].bresp     ),
      .AXI_30_BVALID      (axi3[30].bvalid    ),
      .AXI_31_ACLK        (clk_450            ),
      .AXI_31_ARESET_N    (aresetn_450        ),
      .AXI_31_ARADDR      (axi3[31].araddr    ),
      .AXI_31_ARBURST     (axi3[31].arburst   ),
      .AXI_31_ARID        (axi3[31].arid      ),
      .AXI_31_ARLEN       (axi3[31].arlen     ),
      .AXI_31_ARSIZE      (axi3[31].arsize    ),
      .AXI_31_ARVALID     (axi3[31].arvalid   ),
      .AXI_31_AWADDR      (axi3[31].awaddr    ),
      .AXI_31_AWBURST     (axi3[31].awburst   ),
      .AXI_31_AWID        (axi3[31].awid      ),
      .AXI_31_AWLEN       (axi3[31].awlen     ),
      .AXI_31_AWSIZE      (axi3[31].awsize    ),
      .AXI_31_AWVALID     (axi3[31].awvalid   ),
      .AXI_31_RREADY      (axi3[31].rready    ),
      .AXI_31_BREADY      (axi3[31].bready    ),
      .AXI_31_WDATA       (axi3[31].wdata     ),
      .AXI_31_WLAST       (axi3[31].wlast     ),
      .AXI_31_WSTRB       (axi3[31].wstrb     ),
      .AXI_31_WDATA_PARITY(                   ),
      .AXI_31_WVALID      (axi3[31].wvalid    ),
      .AXI_31_ARREADY     (axi3[31].arready   ),
      .AXI_31_AWREADY     (axi3[31].awready   ),
      .AXI_31_RDATA_PARITY(                   ),
      .AXI_31_RDATA       (axi3[31].rdata     ),
      .AXI_31_RID         (axi3[31].rid       ),
      .AXI_31_RLAST       (axi3[31].rlast     ),
      .AXI_31_RRESP       (axi3[31].rresp     ),
      .AXI_31_RVALID      (axi3[31].rvalid    ),
      .AXI_31_WREADY      (axi3[31].wready    ),
      .AXI_31_BID         (axi3[31].bid       ),
      .AXI_31_BRESP       (axi3[31].bresp     ),
      .AXI_31_BVALID      (axi3[31].bvalid    )
     );

endmodule
